// imem.v 指令存储器模块
module imem(
    input wire [31:0] addr,
    output wire [31:0] inst
);
    // 简单的ROM实现
    reg [31:0] rom [0:255];
    assign inst = rom[addr[9:2]];
    initial begin
        // 测试所有R型指令
        rom[0] = 32'h00500093;  // addi x1, x0, 5      (x1 = 5)
        rom[1] = 32'h00200113;  // addi x2, x0, 2      (x2 = 2, 用于移位测试)
        rom[2] = 32'hffc00193;  // addi x3, x0, -4     (x3 = -4)
        
        // 算术运算测试
        rom[3] = 32'h002081b3;  // add  x3, x1, x2     (x3 = 5 + 2 = 7)
        rom[4] = 32'h40110233;  // sub  x4, x2, x1     (x4 = 2 - 5 = -3)
        
        // 逻辑运算测试
        rom[5] = 32'h0020e2b3;  // or   x5, x1, x2     (x5 = 5 | 2 = 7)
        rom[6] = 32'h0020f333;  // and  x6, x1, x2     (x6 = 5 & 2 = 0)
        rom[7] = 32'h0020c3b3;  // xor  x7, x1, x2     (x7 = 5 ^ 2 = 7)
        
        // 移位运算测试 (x2=2)
        rom[8] = 32'h00209433;  // sll  x8, x1, x2     (x8 = 5 << 2 = 20)
        rom[9] = 32'h0020d4b3;  // srl  x9, x1, x2     (x9 = 5 >> 2 = 1) 
        rom[10] = 32'h4020d533; // sra  x10, x1, x2    (x10 = 5 >>> 2 = 1)
        
        // 比较运算测试
        rom[11] = 32'h0020a5b3; // slt  x11, x1, x2    (x11 = (5 < 2) = 0)
        rom[12] = 32'h0020b633; // sltu x12, x1, x2    (x12 = (5 < 2) = 0)
        
        // 内存操作
        rom[13] = 32'h00302023; // sw   x3, 0(x0)      (存储x3到地址0)
        rom[14] = 32'h00002683; // lw   x13, 0(x0)     (从地址0加载到x13)
        
        // 分支测试
        rom[15] = 32'h00d30463; // beq  x6, x13, +8    (如果x6 == x13则跳转)
        rom[16] = 32'h06300713; // addi x14, x0, 99    (跳过这条)
        rom[17] = 32'h02a00713; // addi x14, x0, 42    (执行这条)
        
        // 死循环
        rom[18] = 32'h00000063; // beq x0, x0, 0       (死循环)
    end
endmodule 