// fibonacci_imem.v - 斐波那契数列计算专用指令存储器
module fibonacci_imem(
    input wire [31:0] addr,
    output wire [31:0] inst
);
    // 简单的ROM实现
    reg [31:0] rom [0:255];
    assign inst = rom[addr[9:2]];
    
    integer i;
    
    initial begin
        // 斐波那契数列计算程序
        // 寄存器分配：
        // x1: fib(n-2) - 第一个斐波那契数
        // x2: fib(n-1) - 第二个斐波那契数  
        // x3: fib(n)   - 当前斐波那契数
        // x4: 计数器 n
        // x5: 最大计数值 (计算到第几个数)
        // x6: 临时寄存器
        // x10: 存储地址计数器
        // x31: 存储基地址
        
        // 初始化
        rom[0] = 32'h00100093;  // addi x1, x0, 1      (fib(0) = 1, 初始化第一个数)
        rom[1] = 32'h00100113;  // addi x2, x0, 1      (fib(1) = 1, 初始化第二个数)  
        rom[2] = 32'h00200213;  // addi x4, x0, 2      (n = 2, 计数器从2开始)
        rom[3] = 32'h00a00293;  // addi x5, x0, 10     (计算到第10个斐波那契数)
        rom[4] = 32'h00000513;  // addi x10, x0, 0     (存储地址计数器 = 0)
        
        // 存储前两个斐波那契数
        rom[5] = 32'h00102023;  // sw x1, 0(x0)        (存储fib(0)=1到地址0)
        rom[6] = 32'h00202223;  // sw x2, 4(x0)        (存储fib(1)=1到地址4)
        rom[7] = 32'h00800513;  // addi x10, x0, 8     (下一个存储地址=8)
        
        // 主循环：计算 fib(n) = fib(n-1) + fib(n-2)
        // 循环入口 (地址 8*4 = 32, 即指令rom[8])
        rom[8] = 32'h002081b3;  // add x3, x1, x2      (x3 = fib(n-2) + fib(n-1))
        
        // 存储当前斐波那契数到内存
        rom[9] = 32'h00352023;  // sw x3, 0(x10)       (存储fib(n)到当前地址)
        
        // 更新斐波那契数：fib(n-2) = fib(n-1), fib(n-1) = fib(n)
        rom[10] = 32'h00010093; // addi x1, x2, 0      (x1 = x2, fib(n-2) = fib(n-1))
        rom[11] = 32'h00018113; // addi x2, x3, 0      (x2 = x3, fib(n-1) = fib(n))
        
        // 递增计数器和地址
        rom[12] = 32'h00120213; // addi x4, x4, 1      (n = n + 1)
        rom[13] = 32'h00450513; // addi x10, x10, 4    (下一个存储地址 += 4)
        
        // 检查是否完成计算
        rom[14] = 32'hfe5244e3; // blt x4, x5, -24     (如果 n < 10，跳转回循环开始rom[8])
        
        // 计算完成，展示结果
        // 依次从内存加载斐波那契数到寄存器x15-x24
        rom[15] = 32'h00002783; // lw x15, 0(x0)       (加载fib(0))
        rom[16] = 32'h00402803; // lw x16, 4(x0)       (加载fib(1))
        rom[17] = 32'h00802883; // lw x17, 8(x0)       (加载fib(2))
        rom[18] = 32'h00c02903; // lw x18, 12(x0)      (加载fib(3))
        rom[19] = 32'h01002983; // lw x19, 16(x0)      (加载fib(4))
        rom[20] = 32'h01402a03; // lw x20, 20(x0)      (加载fib(5))
        rom[21] = 32'h01802a83; // lw x21, 24(x0)      (加载fib(6))
        rom[22] = 32'h01c02b03; // lw x22, 28(x0)      (加载fib(7))
        rom[23] = 32'h02002b83; // lw x23, 32(x0)      (加载fib(8))
        rom[24] = 32'h02402c03; // lw x24, 36(x0)      (加载fib(9))
        
        // 计算结束，进入无限循环
        rom[25] = 32'h00000063; // beq x0, x0, 0       (死循环)
        
        // 剩余位置初始化为NOP
        for (i = 26; i < 256; i = i + 1) begin
            rom[i] = 32'h00000013; // addi x0, x0, 0 (NOP)
        end
    end
endmodule
